module top(
  output wire red_light
);
  assign red_light = 1'b1;       // tie the pin high
endmodule


// red_light
// yellow_light
// green_light