module top(
  output wire red_led
);
  assign red_led = 1'b1;       // tie the pin high
endmodule